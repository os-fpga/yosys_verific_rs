/nfs_scratch/zafar/Castor_V2/DV/unit_level/bram_verif_uvm_env/src/rtl/bram.svh