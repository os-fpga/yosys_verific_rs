`include "/nfs_scratch/scratch/FV/ayyaz/BRAM_TEST1024x2/SIM/bram_rtl.sv"                             
`include "/nfs_scratch/zafar/Castor_V2/DV/unit_level/bram_verif_uvm_env/src/rtl/PLMUX.sv"     
//`include "/nfs_scratch/zafar/Castor_V2/DV/unit_level/bram_verif_uvm_env/src/rtl/ql_clkmux_net.v"  
`include "/nfs_scratch/zafar/Castor_V2/DV/unit_level/bram_verif_uvm_env/src/rtl/sram1024x18.sv"  
`include "/nfs_scratch/zafar/Castor_V2/DV/unit_level/bram_verif_uvm_env/src/rtl/TDP36K.sv"      
`include "/nfs_scratch/zafar/Castor_V2/DV/unit_level/bram_verif_uvm_env/src/rtl/ufifo_ctl.sv"
//`include "/nfs_scratch/zafar/Castor_V2/DV/unit_level/bram_verif_uvm_env/src/rtl/dti_dp_tm16ffcll_1024x18_t8bw2x_m_hc.v"  
//`include "/nfs_scratch/zafar/Castor_V2/DV/unit_level/bram_verif_uvm_env/src/rtl/plmux_top.v"  
`include "/nfs_scratch/zafar/Castor_V2/DV/unit_level/bram_verif_uvm_env/src/rtl/ql_clkmux.v"      
`include "/nfs_scratch/zafar/Castor_V2/DV/unit_level/bram_verif_uvm_env/src/rtl/TDP18K_FIFO.sv"  
`include "/nfs_scratch/zafar/Castor_V2/DV/unit_level/bram_verif_uvm_env/src/rtl/TDP36K_top.sv"
`include "/nfs_scratch/zafar/Castor_V2/DV/unit_level/bram_verif_uvm_env/src/rtl/dti_dp_tm16ffcll_1024x18_t8bw2x_m_hc.v"
//`include "/nfs_scratch/zafar/Castor_V2/DV/unit_level/bram_verif_uvm_env/src/tcbn16ffcllbwp7d5t16p96cpd.v"
//`include "/nfs_scratch/zafar/Castor_V2/DV/unit_level/bram_verif_uvm_env/src/tcbn16ffcllbwp7d5t16p96cpdlvt.v"

