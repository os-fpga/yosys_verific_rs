
(* blackbox *)
module gclkbuff (
    input  A,
    output Z
);

  assign Z = A;

endmodule

