/* Verilog Model Created from SCS Schematic quad_buff.sch 
   Jun 05, 2007 13:39 */

`timescale 1ns/1ns   

module quad_buff( buffer_in , buffer_out );
input buffer_in;
output buffer_out;

assign buffer_out = buffer_in;
endmodule // logic_cell_macro


