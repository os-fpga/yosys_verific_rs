/////////////////////////////////////////
//  Functionality: feedthrough path
//  Author:        George Chen
////////////////////////////////////////
// `timescale 1ns / 1ps


module ft( din, dout);

  input din;
  output dout;

  assign dout = din ;
   
endmodule
