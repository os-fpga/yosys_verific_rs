`ifdef r1024x9_1024x9
`else
`define r1024x9_1024x9
/************************************************************************
** File : r1024x9_1024x9.v
** Design Date: April 11 2006
** Creation Date: Wed Feb 12 10:28:19 2014

** Created By SpDE Version: SpDE 2013.2 Release Build
** Author: QuickLogic Corporation,
** Copyright (C) 1998, Customers of QuickLogic may copy and modify this
** file for use in designing QuickLogic devices only.
** Description : This file is autogenerated RTL code that describes the
** top level design for RAM using QuickLogic's
** RAM block resources.
************************************************************************/
module r1024x9_1024x9 (WA,RA,WD,WD_SEL,RD_SEL,WClk,RClk,WClk_En,RClk_En,WEN,RD);


input [9:0] WA;
input [9:0] RA;
input WD_SEL,RD_SEL;
input WClk,RClk;
input WClk_En,RClk_En;
input [0:0] WEN;
input [8:0] WD;
output [8:0] RD;

reg [8:0] RAM9bit;
wire WEN01;
wire V_clk;

assign V_clk = WClk | RClk;
assign WEN01 = WEN | WD_SEL;
assign RD = ((RD_SEL == 1'b1 ) && (RClk_En == 1'b1)) ? RAM9bit : 16'b0;

always @(posedge V_clk)
begin
	if ((WD_SEL == 1'b1 ) && (WClk_En == 1'b1) && (WEN01 == 1'b1 ))
	RAM9bit <= {WA,RA,WD_SEL,RD_SEL} ^ WD;
end

endmodule
`endif


//module RAM_RW(WA,RA,WD,WD_SEL,RD_SEL,WClk,RClk,WClk_En,RClk_En,WEN,RD); 
